module memory(clk,reset,data_in,n_valid,valid_state,pathVec,ifFinal);
input clk;
input reset;
input [9:0] data_in;
input n_valid;

output [9:0] valid_state;
output [31:0] pathVec;
output ifFinal;

wire clk;
wire reset;
wire [9:0] data_in;
wire n_valid;

reg [9:0] valid_state;
reg [31:0] pathVec;
reg ifFinal;

reg [40:0] mem_in[0:1023];

always@(posedge clk)
begin
	if(reset == 1)
	begin
		valid_state <= 0;
		pathVec     <= 32'b11111111111111111111111111111111;
	   	ifFinal     <= 0;	
   mem_in[8'b00000001] <= { 1'b0, 8'b00000001 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000010] <= { 1'b0, 8'b00000010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00100101] <= { 1'b0, 8'b00100101 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00101100] <= { 1'b0, 8'b00101100 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000010] <= { 1'b0, 8'b00000010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000010] <= { 1'b0, 8'b00000010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000010] <= { 1'b0, 8'b00000010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000010] <= { 1'b0, 8'b00000010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b01100100] <= { 1'b0, 8'b01100100 ,32'b11111111111111111111111111111111 };
   mem_in[8'b01101011] <= { 1'b0, 8'b01101011 ,32'b11111111111111111111111111111111 };
   mem_in[8'b01110010] <= { 1'b0, 8'b01110010 ,32'b11111111111111111111111111111111 };
   mem_in[8'b01111001] <= { 1'b0, 8'b01111001 ,32'b11111111111111111111111111111111 };
   mem_in[8'b10001110] <= { 1'b0, 8'b10001110 ,32'b11111111111111111111111111111111 };
   mem_in[8'b10010101] <= { 1'b0, 8'b10010101 ,32'b11111111111111111111111111111111 };
   mem_in[8'b00000011] <= { 1'b0, 8'b00000011 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00000100] <= { 1'b0, 8'b00000100 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00000101] <= { 1'b0, 8'b00000101 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00000110] <= { 1'b0, 8'b00000110 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00000111] <= { 1'b0, 8'b00000111 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00001000] <= { 1'b1, 8'b00001000 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00011101] <= { 1'b1, 8'b00011101 ,32'b00000000000000000000001000001001 };
   mem_in[8'b00001010] <= { 1'b0, 8'b00001010 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00001011] <= { 1'b0, 8'b00001011 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00001100] <= { 1'b0, 8'b00001100 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00001101] <= { 1'b0, 8'b00001101 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00001110] <= { 1'b0, 8'b00001110 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00001111] <= { 1'b1, 8'b00001111 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00010110] <= { 1'b1, 8'b00010110 ,32'b00000000000000000010110000010110 };
   mem_in[8'b00100100] <= { 1'b1, 8'b00100100 ,32'b00000000000000000010110000010000 };
   mem_in[8'b00100110] <= { 1'b0, 8'b00100110 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00100111] <= { 1'b0, 8'b00100111 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00101000] <= { 1'b0, 8'b00101000 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00101001] <= { 1'b0, 8'b00101001 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00101010] <= { 1'b0, 8'b00101010 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00101011] <= { 1'b1, 8'b00101011 ,32'b00000000000000000000000000100000 };
   mem_in[8'b00101101] <= { 1'b0, 8'b00101101 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00101110] <= { 1'b0, 8'b00101110 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00101111] <= { 1'b0, 8'b00101111 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00110000] <= { 1'b0, 8'b00110000 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00110001] <= { 1'b0, 8'b00110001 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00110010] <= { 1'b1, 8'b00110010 ,32'b00000000000000000000000001000000 };
   mem_in[8'b00110100] <= { 1'b0, 8'b00110100 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00110101] <= { 1'b0, 8'b00110101 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00110110] <= { 1'b0, 8'b00110110 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00110111] <= { 1'b0, 8'b00110111 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00111000] <= { 1'b0, 8'b00111000 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00111001] <= { 1'b1, 8'b00111001 ,32'b00000000000000000000000010000000 };
   mem_in[8'b00111011] <= { 1'b0, 8'b00111011 ,32'b00000000000000000000000100000000 };
   mem_in[8'b00111100] <= { 1'b0, 8'b00111100 ,32'b00000000000000000000000100000000 };
   mem_in[8'b00111101] <= { 1'b0, 8'b00111101 ,32'b00000000000000000000000100000000 };
   mem_in[8'b00111110] <= { 1'b0, 8'b00111110 ,32'b00000000000000000000000100000000 };
   mem_in[8'b00111111] <= { 1'b0, 8'b00111111 ,32'b00000000000000000000000100000000 };
   mem_in[8'b01000000] <= { 1'b1, 8'b01000000 ,32'b00000000000000000000000100000000 };
   mem_in[8'b01010111] <= { 1'b0, 8'b01010111 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01011000] <= { 1'b0, 8'b01011000 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01011001] <= { 1'b0, 8'b01011001 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01011010] <= { 1'b0, 8'b01011010 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01011011] <= { 1'b0, 8'b01011011 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01011100] <= { 1'b1, 8'b01011100 ,32'b00000000000000000001000000000000 };
   mem_in[8'b01100101] <= { 1'b0, 8'b01100101 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01100110] <= { 1'b0, 8'b01100110 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01100111] <= { 1'b0, 8'b01100111 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01101000] <= { 1'b0, 8'b01101000 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01101001] <= { 1'b0, 8'b01101001 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01101010] <= { 1'b1, 8'b01101010 ,32'b00000000000000000100000000000000 };
   mem_in[8'b01101100] <= { 1'b0, 8'b01101100 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01101101] <= { 1'b0, 8'b01101101 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01101110] <= { 1'b0, 8'b01101110 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01101111] <= { 1'b0, 8'b01101111 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01110000] <= { 1'b0, 8'b01110000 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01110001] <= { 1'b1, 8'b01110001 ,32'b00000000000000001000000000000000 };
   mem_in[8'b01110011] <= { 1'b0, 8'b01110011 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01110100] <= { 1'b0, 8'b01110100 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01110101] <= { 1'b0, 8'b01110101 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01110110] <= { 1'b0, 8'b01110110 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01110111] <= { 1'b0, 8'b01110111 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01111000] <= { 1'b1, 8'b01111000 ,32'b00000000000000010000000000000000 };
   mem_in[8'b01111010] <= { 1'b0, 8'b01111010 ,32'b00000000000000100000000000000000 };
   mem_in[8'b01111011] <= { 1'b0, 8'b01111011 ,32'b00000000000000100000000000000000 };
   mem_in[8'b01111100] <= { 1'b0, 8'b01111100 ,32'b00000000000000100000000000000000 };
   mem_in[8'b01111101] <= { 1'b0, 8'b01111101 ,32'b00000000000000100000000000000000 };
   mem_in[8'b01111110] <= { 1'b0, 8'b01111110 ,32'b00000000000000100000000000000000 };
   mem_in[8'b01111111] <= { 1'b1, 8'b01111111 ,32'b00000000000000100000000000000000 };
   mem_in[8'b10000001] <= { 1'b0, 8'b10000001 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10000010] <= { 1'b0, 8'b10000010 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10000011] <= { 1'b0, 8'b10000011 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10000100] <= { 1'b0, 8'b10000100 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10000101] <= { 1'b0, 8'b10000101 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10000110] <= { 1'b1, 8'b10000110 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10001101] <= { 1'b1, 8'b10001101 ,32'b00000000000011000000000000000000 };
   mem_in[8'b10001111] <= { 1'b0, 8'b10001111 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010000] <= { 1'b0, 8'b10010000 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010001] <= { 1'b0, 8'b10010001 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010010] <= { 1'b0, 8'b10010010 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010011] <= { 1'b0, 8'b10010011 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010100] <= { 1'b1, 8'b10010100 ,32'b00000000000100000000000000000000 };
   mem_in[8'b10010110] <= { 1'b0, 8'b10010110 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10010111] <= { 1'b0, 8'b10010111 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10011000] <= { 1'b0, 8'b10011000 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10011001] <= { 1'b0, 8'b10011001 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10011010] <= { 1'b0, 8'b10011010 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10011011] <= { 1'b1, 8'b10011011 ,32'b00000000001000000000000000000000 };
   mem_in[8'b10011101] <= { 1'b0, 8'b10011101 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10011110] <= { 1'b0, 8'b10011110 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10011111] <= { 1'b0, 8'b10011111 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10100000] <= { 1'b0, 8'b10100000 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10100001] <= { 1'b0, 8'b10100001 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10100010] <= { 1'b1, 8'b10100010 ,32'b00000000010000000000000000000000 };
   mem_in[8'b10100100] <= { 1'b0, 8'b10100100 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10100101] <= { 1'b0, 8'b10100101 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10100110] <= { 1'b0, 8'b10100110 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10100111] <= { 1'b0, 8'b10100111 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10101000] <= { 1'b0, 8'b10101000 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10101001] <= { 1'b1, 8'b10101001 ,32'b00000000100000000000000000000000 };
   mem_in[8'b10101011] <= { 1'b0, 8'b10101011 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10101100] <= { 1'b0, 8'b10101100 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10101101] <= { 1'b0, 8'b10101101 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10101110] <= { 1'b0, 8'b10101110 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10101111] <= { 1'b0, 8'b10101111 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10110000] <= { 1'b1, 8'b10110000 ,32'b00000001000000000000000000000000 };
   mem_in[8'b10110010] <= { 1'b0, 8'b10110010 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10110011] <= { 1'b0, 8'b10110011 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10110100] <= { 1'b0, 8'b10110100 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10110101] <= { 1'b0, 8'b10110101 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10110110] <= { 1'b0, 8'b10110110 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10110111] <= { 1'b1, 8'b10110111 ,32'b00000010000000000000000000000000 };
   mem_in[8'b10111001] <= { 1'b0, 8'b10111001 ,32'b00000100000000000000000000000000 };
   mem_in[8'b10111010] <= { 1'b0, 8'b10111010 ,32'b00000100000000000000000000000000 };
   mem_in[8'b10111011] <= { 1'b0, 8'b10111011 ,32'b00000100000000000000000000000000 };
   mem_in[8'b10111100] <= { 1'b0, 8'b10111100 ,32'b00000100000000000000000000000000 };
   mem_in[8'b10111101] <= { 1'b0, 8'b10111101 ,32'b00000100000000000000000000000000 };
   mem_in[8'b10111110] <= { 1'b1, 8'b10111110 ,32'b00000100000000000000000000000000 };
   mem_in[8'b11000000] <= { 1'b0, 8'b11000000 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000001] <= { 1'b0, 8'b11000001 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000010] <= { 1'b0, 8'b11000010 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000011] <= { 1'b0, 8'b11000011 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000100] <= { 1'b0, 8'b11000100 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000101] <= { 1'b1, 8'b11000101 ,32'b00001000000000000000000000000000 };
   mem_in[8'b11000111] <= { 1'b0, 8'b11000111 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001000] <= { 1'b0, 8'b11001000 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001001] <= { 1'b0, 8'b11001001 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001010] <= { 1'b0, 8'b11001010 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001011] <= { 1'b0, 8'b11001011 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001100] <= { 1'b1, 8'b11001100 ,32'b00010000000000000000000000000000 };
   mem_in[8'b11001110] <= { 1'b0, 8'b11001110 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11001111] <= { 1'b0, 8'b11001111 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11010000] <= { 1'b0, 8'b11010000 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11010001] <= { 1'b0, 8'b11010001 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11010010] <= { 1'b0, 8'b11010010 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11010011] <= { 1'b1, 8'b11010011 ,32'b00100000000000000000000000000000 };
   mem_in[8'b11010101] <= { 1'b0, 8'b11010101 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11010110] <= { 1'b0, 8'b11010110 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11010111] <= { 1'b0, 8'b11010111 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11011000] <= { 1'b0, 8'b11011000 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11011001] <= { 1'b0, 8'b11011001 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11011010] <= { 1'b1, 8'b11011010 ,32'b01000000000000000000000000000000 };
   mem_in[8'b11011100] <= { 1'b0, 8'b11011100 ,32'b10000000000000000000000000000000 };
   mem_in[8'b11011101] <= { 1'b0, 8'b11011101 ,32'b10000000000000000000000000000000 };
   mem_in[8'b11011110] <= { 1'b0, 8'b11011110 ,32'b10000000000000000000000000000000 };
   mem_in[8'b11011111] <= { 1'b0, 8'b11011111 ,32'b10000000000000000000000000000000 };
   mem_in[8'b11100000] <= { 1'b0, 8'b11100000 ,32'b10000000000000000000000000000000 };
   mem_in[8'b11100001] <= { 1'b1, 8'b11100001 ,32'b10000000000000000000000000000000 };
   end

   else if(n_valid == 1)
   	begin 
	   valid_state <= 0;
	   pathVec     <= 32'b11111111111111111111111111111111;
	   ifFinal     <= 0;	
	end
  else	
   	begin 
	   valid_state <= mem_in[data_in][39:32];
	   pathVec     <= mem_in[data_in][31:0];
	   ifFinal     <= mem_in[data_in][40];	
	end   
   end
   
   
endmodule   
	   
	   
